//=====================================================================
//  FILES REQUIRED FOR FIFO TESTBENCH
//=====================================================================
//
//  signals.sv        : Contains parameter definitions and I/O signal declarations
//  clk_gen.sv        : Clock generator class for driving the testbench clock
//  reset_gen.sv      : Reset generator class (if separate)
//  condition_test.sv : Contains write/read tasks, functional checks,
//                      and condition-specific test scenarios
//  run.sv            : Main test sequence class that coordinates
//                      reset, stimulus generation, checks, and reporting
//
//=====================================================================

`include "signals.sv"
`include "clk_gen.sv"
`include "reset_gen.sv"      // (Add if you use a separate reset file)
`include "condition_test.sv"
`include "run.sv"